`timescale 1ns/1ps
module fifo_tb();

endmodule